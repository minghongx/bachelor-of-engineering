module entry_indicator (
	input rst_ni,
	input entry_i,
	output entering_last_digit_o
);

endmodule
